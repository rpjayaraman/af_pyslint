class add;
  bit var1;
endclass :add 
